`timescale 1ns / 1ps


module tb_factorial #(parameter DATA_WIDTH = 4);
    reg clk_tb, rst_tb;



endmodule