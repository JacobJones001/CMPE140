module factorial #(parameter DATA_WIDTH = 32)(
    input rst, clk,
    input Go,
    input [DATA_WIDTH-1:0] n,
    output Done, Error,
    output [DATA_WIDTH-1:0] product
);





endmodule