module controlunit (
        input  wire [5:0]  opcode,
        input  wire [5:0]  funct,
        output wire        branch,
        output wire        jump,
        output wire        reg_dst,
        output wire        we_reg,
        output wire        alu_src,
        output wire        we_dm,
        output wire        dm2reg,
        output wire        hilo_sel,
        output wire        alu_out_sel,
        output wire        we_hilo,
        output wire [2:0]  alu_ctrl
    );
    
    wire [1:0] alu_op;
    // wire hilo_sel;
    // wire dm2reg_0;
    // assign dm2reg = {hilo_sel, dm2reg_0};

    maindec md (
        .opcode         (opcode),
        .branch         (branch),
        .jump           (jump),
        .reg_dst        (reg_dst),
        .we_reg         (we_reg),
        .alu_src        (alu_src),
        .we_dm          (we_dm),
        .dm2reg         (dm2reg),
        .alu_op         (alu_op)
    );

    auxdec ad (
        .alu_op         (alu_op),
        .funct          (funct),
        .alu_ctrl       (alu_ctrl),
        .hilo_sel       (hilo_sel),
        .alu_out_sel    (alu_out_sel)
    );

endmodule